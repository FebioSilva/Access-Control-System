library ieee;
use ieee.std_logic_1164.all;

entity SLCDC_tb is
	end SLCDC_tb;
	
architecture behavioral of SLCDC_tb is

component SLCDC is
  port(
	 SDX: in std_logic;
   SCLK: in std_logic;
   SS: in std_logic;
   rst : in std_logic;
	clk : in std_logic;
	
	Wrl: out std_logic;
	Dout: out std_logic_vector(4 downto 0)
    );
end component SLCDC;

constant MCLK_PERIOD : time :=20ns;
constant	MCLK_HALF_PERIOD : time :=MCLK_PERIOD/2;

signal SDX_tb, SS_tb,SCLK_tb,clk_tb,rst_tb,Wrl_tb : std_logic;
signal Dout_tb : std_logic_vector(4 downto 0);

begin

UUT: SLCDC port map(SDX => SDX_tb,
						  SS => SS_tb,
                    clk => clk_tb,
                    rst => rst_tb,
                    Wrl => Wrl_tb,
						  SCLK => SCLK_tb,
						  Dout => Dout_tb
						  );
clk_gen : process
begin
	clk_tb <= '0';
	wait for MCLK_HALF_PERIOD/2;
	clk_tb <= '1';
	wait for MCLK_HALF_PERIOD/2;
end process;

clk_gen2 : process
begin
	SCLK_tb <= '0';
	wait for MCLK_HALF_PERIOD;
	SCLK_tb <= '1';
	wait for MCLK_HALF_PERIOD;
end process;

stimulus: process
begin
    SDX_tb <= '1';
	 SS_tb <= '1';
	 rst_tb <= '1';
	wait for MCLK_PERIOD;
	
	  rst_tb <= '0';
	  SS_tb <='0';	
	wait for 5*MCLK_PERIOD;

	  SS_tb <= '1';
	wait for 4*MCLK_PERIOD;
	
	wait;
end process;
end behavioral;

		