library ieee;
use ieee.std_logic_1164.all;

entity KeyDecoder_tb is
	end KeyDecoder_tb;
	
architecture behavioral of KeyDecoder_tb is

component KeyDecoder is
port(
	Kack : in std_logic;
	CLK : in std_logic;
	Rst : in std_logic;
	Ln1,Ln2,Ln3, Ln4: in std_logic;
	
	Col1,Col2,Col3: out std_logic;
	Kval : out std_logic;
	K : out std_logic_vector(3 downto 0)
	);
end component KeyDecoder;

constant MCLK_PERIOD : time :=20ns;
constant	MCLK_HALF_PERIOD : time :=MCLK_PERIOD/2;

signal Kack_tb,CLK_tb,Rst_tb,Ln1_tb,Ln2_tb,Ln3_tb,Ln4_tb,Col1_tb,Col2_tb,Col3_tb,Kval_tb : std_logic;
signal K_tb : std_logic_vector(3 downto 0);
begin

UUT: KeyDecoder port map(Kack => Kack_tb, 
							 CLK => CLK_tb, 
							 Rst => Rst_tb, 
							 Ln1 => Ln1_tb,
							 Ln2 => Ln2_tb,
							 Ln3 => Ln3_tb, 
							 Ln4 => Ln4_tb,
							 Col1 => Col1_tb,
							 Col2 => Col2_tb,
							 Col3 => Col3_tb,
							 Kval => Kval_tb,
							 K => K_tb
							 );
clk_gen : process
begin
	clk_tb <= '0';
	wait for MCLK_HALF_PERIOD;
	clk_tb <= '1';
	wait for MCLK_HALF_PERIOD;
end process;

stimulus: process
begin
	Kack_tb <= '0';
	Rst_tb <= '1';
	Ln1_tb <='1';
	Ln2_tb <='1';
	Ln3_tb <='1';
	Ln4_tb <='1';
	wait for MCLK_PERIOD;
	
	
	Rst_tb <='0';
	Kack_tb <='1';
	wait for MCLK_PERIOD;
	
	Ln1_tb <='0';
	wait for 3*MCLK_PERIOD;
	
	Kack_tb <= '0';
	Ln1_tb <='1';
	wait for MCLK_PERIOD;
	
	Kack_tb <= '1';
	Ln2_tb <= '0';
	wait for 3*MCLK_PERIOD;
	
	Kack_tb <= '0';
	Ln2_tb <='1';
	wait for 2*MCLK_PERIOD;
	
	Kack_tb <= '1';
	Ln3_tb <='0';
	wait for 3*MCLK_PERIOD;
	
	Kack_tb <= '0';
	Ln3_tb <='1';
	wait for MCLK_PERIOD;	
	wait;
end process;
end behavioral;

		