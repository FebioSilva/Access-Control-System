library ieee;
use ieee.std_logic_1164.all;

entity MAC_tb is
	end MAC_tb;
	
architecture behavioral of MAC_tb is

component MAC is
	port(
	putget: in std_logic;
	incPut: in std_logic;
	incGet: in std_logic;
	clk: in std_logic;
	reset: in std_logic;
	
	full: out std_logic;
	empty: out std_logic;
	Aout: out std_logic_vector(2 downto 0)
	);
end component MAC;

constant MCLK_PERIOD : time :=20ns;
constant	MCLK_HALF_PERIOD : time :=MCLK_PERIOD/2;

signal full_tb, empty_tb, reset_tb, clk_tb, putget_tb, incGet_tb, incPut_tb : std_logic;
signal Aout_tb: std_logic_vector(2 downto 0);

begin

UUT: MAC port map(full => full_tb, empty => empty_tb, reset => reset_tb, clk => clk_tb,
										  incGet => incGet_tb, incPut => incPut_tb, putget => putget_tb, Aout => Aout_tb
										  );
clk_gen : process
begin
	clk_tb <= '0';
	wait for MCLK_HALF_PERIOD;
	clk_tb <= '1';
	wait for MCLK_HALF_PERIOD;
end process;


stimulus: process
begin
	putget_tb <= '0';
	incPut_tb <= '0';
	incGet_tb <= '0';
	reset_tb <='1';
	wait for MCLK_PERIOD;
	
	putget_tb <= '1';
	incPut_tb <= '1';
	reset_tb <='0';
	wait for 8*MCLK_PERIOD;
	
	putget_tb <= '0';
	incPut_tb <= '0';
	wait for MCLK_PERIOD;
	
	
	incGet_tb <= '1';
	wait for 8*MCLK_PERIOD;
	
	incGet_tb <= '0';
	wait for MCLK_PERIOD;
	
	wait for MCLK_PERIOD;
	wait;
end process;
end behavioral;

		