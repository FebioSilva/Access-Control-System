LIBRARY IEEE;
use IEEE.std_logic_1164.all;

entity PEnc4 is 
	port
	(
	A : in std_logic_vector(3 downto 0);--I
	R : out std_logic_vector(1 downto 0);--O
	V : out std_logic--V
	);
end Penc4;

architecture structural of Penc4 is begin
	R(0) <= (A(1) AND NOT A(2)) OR A(3); --A(1) and (not A(2)) or A(3); Se quisermos modificar para less significant input
	R(1) <= A(2) OR A(3);
	V <= A(0) OR A(1) OR A(2) OR A(3);
	
end structural; 